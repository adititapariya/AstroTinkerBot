module AND_GATE (
    input a,b,          // defining inputs A and B of AND gate
    output out          // defining output of AND gate
);

assign out = a & b;     // Logic implementation

endmodule
